module norgate(a,b,c) ;
input a,b;
output c;
nor a1(c,a,b);

    
endmodule