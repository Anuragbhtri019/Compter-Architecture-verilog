module nandgate ( a,b,c) ;
input a,b;
output c;
nand n1(c,a,b);   
endmodule