 module orgate(a,b,c);
 input a,b;
 output c;
 or a1(c,a,b);
endmodule