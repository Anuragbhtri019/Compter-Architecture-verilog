module xnorgate(a,b,c);
input a,b;
output c;
xnor a1(c,a,b);
endmodule