module xorgate(a,b,c);
input a,b;
output  c;
xor a1(c,a,b);
endmodule