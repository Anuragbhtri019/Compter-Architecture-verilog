module andgate(a,b,c);
input a,b;
output c;
and a1(c,a,b);
endmodule