module notgate(a,c);
input a;
output c;
not a1(c,a);
endmodule;